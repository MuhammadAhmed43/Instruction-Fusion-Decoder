module core #(
    parameter FUSION_ENABLE = 1
)(
    input wire clk,
    input wire rst,
    input wire data_mem_valid,
    input wire instruc_mem_valid,
    input wire [31:0] instruction,
    input wire [31:0] load_data_in,

    output wire load_signal,
    output wire instruction_mem_we_re,
    output wire instruction_mem_request,
    output wire data_mem_we_re,
    output wire data_mem_request,
    output wire [3:0]  mask_singal,
    output wire [3:0]  instruc_mask_singal,
    output wire [31:0] store_data_out,
    output wire [31:0] alu_out_address,
    output wire [31:0] pc_address
    );

    wire [31:0] instruc_data_out;
    wire [31:0] pre_address_pc;
    wire [31:0] instruction_fetch , instruction_decode , instruction_execute;
    wire [31:0] instruction_memstage , instruction_wb;
    wire [31:0] pre_pc_addr_fetch , pre_pc_addr_decode , pre_pc_addr_execute;
    wire [31:0] pre_pc_addr_memstage , pre_pc_addr_wb;
    wire load_decode , load_execute , load_memstage;
    wire store_decode , store_execute , store_memstage;
    wire jalr_decode;
    wire next_sel_decode , next_sel_execute;
    wire reg_write_decode , reg_write_execute , reg_write_memstage;
    wire branch_result_decode , branch_result_execute;
    wire [3:0]  mask;
    wire [3:0]  alu_control_decode , alu_control_execute;
    wire [1:0]  mem_to_reg_decode , mem_to_reg_execute;
    wire [1:0]  mem_to_reg_memstage , mem_to_reg_wb;
    wire [4:0]  rs1_decode , rs1_execute;
    wire [4:0]  rs2_decode , rs2_execute;
    wire [4:0]  rd_memstage;
    wire [31:0] op_b_decode , op_b_execute , op_b_memstage;
    wire [31:0] opa_mux_out_decode , opa_mux_out_execute;
    wire [31:0] opb_mux_out_decode , opb_mux_out_execute;
    wire [31:0] alu_res_out_execute , alu_res_out_memstage;
    wire [31:0] alu_res_out_wb;
    wire [31:0] next_sel_address_execute , next_sel_address_memstage;
    wire [31:0] next_sel_address_wb;
    wire [31:0] wrap_load_memstage , wrap_load_wb;
    wire [31:0] rd_wb_data;
    wire [31:0] alu_in_a , alu_in_b;
    wire operand_a_decode, operand_b_decode;
    wire operand_a_execute, operand_b_execute;
    
    // FUSION SIGNALS
    wire fuse_flag_raw;
    wire fuse_flag;
    wire [1:0] fuse_type;
    wire [31:0] fused_inst;
    wire hazard_stall;

    // Apply fusion only when enabled
    assign fuse_flag = fuse_flag_raw & FUSION_ENABLE;
    
    // IMPORTANT: Load+ALU fusion (fuse_type=11) should NOT skip the second instruction!
    // Load+ALU fusion works by forwarding loaded data, both instructions still execute.
    // Only LUI+ADDI (01) and AUIPC+JALR (10) skip the second instruction.
    wire fuse_flag_skip = fuse_flag && (fuse_type != 2'b11);

    // ==========================================================================
    // HAZARD DETECTION (Artificial Stalls for Baseline Comparison)
    // ==========================================================================
    // When Fusion is DISABLED, we enforce stalls on RAW hazards for specific
    // patterns. This simulates a processor without full forwarding for these
    // cases, allowing Fusion to demonstrate speedup by avoiding the stall.
    // ==========================================================================
    
    // LUI -> ADDI hazard (for LUI+ADDI fusion)
    wire lui_addi_hazard = (instruction_execute[6:0] == 7'b0110111) && // LUI in Ex
                           (instruction_decode[6:0] == 7'b0010011) &&  // ADDI in Dec
                           (instruction_execute[11:7] == instruction_decode[19:15]) && // rd == rs1
                           (instruction_execute[11:7] != 0);
    
    // AUIPC -> JALR hazard (for AUIPC+JALR fusion)
    wire auipc_jalr_hazard = (instruction_execute[6:0] == 7'b0010111) && // AUIPC in Ex
                              (instruction_decode[6:0] == 7'b1100111) && // JALR in Dec
                              (instruction_execute[11:7] == instruction_decode[19:15]) && // rd == rs1
                              (instruction_execute[11:7] != 0);
    
    // LOAD -> ALU hazard (for LOAD+ALU fusion)
    wire load_alu_hazard_rs1 = (instruction_execute[6:0] == 7'b0000011) && // Load in Ex
                                ((instruction_decode[6:0] == 7'b0110011) ||  // R-type in Dec
                                 (instruction_decode[6:0] == 7'b0010011)) && // I-type in Dec
                                (instruction_execute[11:7] == instruction_decode[19:15]) && // rd == rs1
                                (instruction_execute[11:7] != 0);
    
    wire load_alu_hazard_rs2 = (instruction_execute[6:0] == 7'b0000011) && // Load in Ex
                                (instruction_decode[6:0] == 7'b0110011) &&  // R-type only
                                (instruction_execute[11:7] == instruction_decode[24:20]) && // rd == rs2
                                (instruction_execute[11:7] != 0);
    
    wire load_alu_hazard = load_alu_hazard_rs1 | load_alu_hazard_rs2;

    // Combined hazard stall (only when fusion is disabled)
    // When fusion is ENABLED, Load+ALU patterns are handled by forwarding loaded data
    assign hazard_stall = (!FUSION_ENABLE) && (lui_addi_hazard | auipc_jalr_hazard | load_alu_hazard);

    //FETCH STAGE
    fetch u_fetchstage(
        .clk(clk),
        .rst(rst),
        .load(load_decode | hazard_stall), // Stall Fetch
        .jalr(jalr_execute),
        .next_sel(next_sel_execute),
        .branch_reselt(branch_result_execute),
        .fuse_skip(fuse_flag_skip),
        .next_address(alu_res_out_execute),
        .instruction_fetch(instruction),
        .instruction(instruction_fetch),
        .address_in(0),
        .valid(data_mem_valid),
        .mask(instruc_mask_singal),
        .we_re(instruction_mem_we_re),
        .request(instruction_mem_request),
        .pre_address_pc(pre_pc_addr_fetch),
        .address_out(pc_address)
    );

    //FETCH STAGE PIPELINE
    fetch_pipe u_fetchpipeline(
        .clk(clk),
        .rst(rst),
        .pre_address_pc(pre_pc_addr_fetch),
        .instruction_fetch(instruction_fetch),
        .pre_address_out(pre_pc_addr_decode),
        .instruction(instruction_decode),
        .next_select(next_sel_decode),
        .branch_result(branch_result_decode),
        .jalr(jalr_decode),
        .load(load_decode | hazard_stall), // Stall Fetch Pipe
        .fuse_flush(fuse_flag_skip)
    );

    // FUSION DECODER
    fusion_decoder u_fusion_decoder(
        .inst1(instruction_decode),
        .inst2(instruction_fetch),
        .fuse_flag(fuse_flag_raw),
        .fuse_type(fuse_type),
        .fused_inst(fused_inst)
    );

    //DECODE STAGE
    decode u_decodestage(
        .clk(clk),
        .rst(rst),
        .valid(data_mem_valid),
        .load_control_signal(load_execute),
        .reg_write_en_in(reg_write_wb),
        .instruction(fuse_flag ? fused_inst : instruction_decode),
        .pc_address(pre_pc_addr_decode),
        .rd_wb_data(rd_wb_data),
        .rs1(rs1_decode),
        .rs2(rs2_decode),
        .load(load_decode),
        .store(store_decode),
        .jalr(jalr_decode),
        .next_sel(next_sel_decode),
        .reg_write_en_out(reg_write_decode),
        .mem_to_reg(mem_to_reg_decode),
        .branch_result(branch_result_decode),
        .opb_data(op_b_decode),
        .instruction_rd(instruction_wb),
        .alu_control(alu_control_decode),
        .opa_mux_out(opa_mux_out_decode),
        .opb_mux_out(opb_mux_out_decode),
        .operand_a_out(operand_a_decode),
        .operand_b_out(operand_b_decode),
        
        // Forwarding Wiring
        .alu_result_execute(alu_res_out_execute),
        .rd_execute(instruction_execute[11:7]),
        .reg_write_execute(reg_write_execute),
        .alu_result_mem(alu_res_out_memstage),
        .rd_mem(rd_memstage),
        .reg_write_mem(reg_write_memstage)
    );

    //DECODE STAGE PIPELINE
    decode_pipe u_decodepipeline(
        .clk(clk),
        .rst(rst),
        .flush(hazard_stall), // Flush Execute (Insert Bubble)
        .load_in(load_decode),
        .store_in(store_decode),
        .jalr_in(jalr_decode),
        .next_sel_in(next_sel_decode),
        .mem_to_reg_in(mem_to_reg_decode),
        .branch_result_in(branch_result_decode),
        .opb_data_in(op_b_decode),
        .alu_control_in(alu_control_decode),
        .opa_mux_in(opa_mux_out_decode),
        .opb_mux_in(opb_mux_out_decode),
        .pre_address_in(pre_pc_addr_decode),
        .instruction_in(instruction_decode),
        .reg_write_in(reg_write_decode),
        .rs1_in(rs1_decode),
        .rs2_in(rs2_decode),
        .operand_a_in(operand_a_decode),
        .operand_b_in(operand_b_decode),
        .reg_write_out(reg_write_execute),
        .jalr_out(jalr_execute),
        .load(load_execute),
        .store(store_execute),
        .next_sel(next_sel_execute),
        .mem_to_reg(mem_to_reg_execute),
        .branch_result(branch_result_execute),
        .opb_data_out(op_b_execute),
        .alu_control(alu_control_execute),
        .opa_mux_out(opa_mux_out_execute),
        .opb_mux_out(opb_mux_out_execute),
        .pre_address_out(pre_pc_addr_execute),
        .instruction_out(instruction_execute),
        .rs1_out(rs1_execute),
        .rs2_out(rs2_execute),
        .operand_a_out(operand_a_execute),
        .operand_b_out(operand_b_execute)
    );

    // Detect if instruction in Memory stage is a Load (opcode 0000011)
    wire load_in_memstage = (instruction_memstage[6:0] == 7'b0000011);
    
    // Select correct data from Memory stage: loaded data for Loads, ALU result otherwise
    wire [31:0] mem_forward_data = load_in_memstage ? wrap_load_memstage : alu_res_out_memstage;

    // Forwarding logic with MEM and WB stages
    // For Load instructions in MEM stage, forward the loaded data (wrap_load_memstage)
    // For other instructions in MEM stage, forward the ALU result (alu_res_out_memstage)
    assign alu_in_a = (!operand_a_execute && rs1_execute == rd_memstage && reg_write_memstage && rd_memstage != 0) ? mem_forward_data : 
                      (!operand_a_execute && rs1_execute == instruction_wb[11:7] && reg_write_wb && instruction_wb[11:7] != 0) ? rd_wb_data :
                      opa_mux_out_execute;

    assign alu_in_b = (!operand_b_execute && rs2_execute == rd_memstage && reg_write_memstage && rd_memstage != 0) ? mem_forward_data :
                      (!operand_b_execute && rs2_execute == instruction_wb[11:7] && reg_write_wb && instruction_wb[11:7] != 0) ? rd_wb_data :
                      opb_mux_out_execute;

    //EXECUTE STAGE
    execute u_executestage(
        .a_i(alu_in_a),
        .b_i(alu_in_b),
        .pc_address(pre_pc_addr_execute),
        .alu_control(alu_control_execute),
        .alu_res_out(alu_res_out_execute),
        .next_sel_address(next_sel_address_execute)
    );

    //EXECUTE STAGE PIPELINE
    execute_pipe u_executepipeline(
        .clk(clk),
        .rst(rst),
        .load_in(load_execute),
        .store_in(store_execute),
        .opb_datain(op_b_execute),
        .alu_res(alu_res_out_execute),
        .mem_reg_in(mem_to_reg_execute),
        .next_sel_addr(next_sel_address_execute),
        .pre_address_in(pre_pc_addr_execute),
        .instruction_in(instruction_execute),
        .reg_write_in(reg_write_execute),
        .reg_write_out(reg_write_memstage),
        .load_out(load_memstage),
        .store_out(store_memstage),
        .opb_dataout(op_b_memstage),
        .alu_res_out(alu_res_out_memstage),
        .mem_reg_out(mem_to_reg_memstage),
        .next_sel_address(next_sel_address_memstage),
        .pre_address_out(pre_pc_addr_memstage),
        .instruction_out(instruction_memstage)
    );

    //MEMORY STAGE
    memory_stage u_memorystage(
        .rst(rst),
        .load(load_memstage),
        .store(store_memstage),
        .op_b(op_b_memstage),
        .instruction(instruction_memstage),
        .alu_out_address(alu_res_out_memstage),
        .wrap_load_in(load_data_in),
        .mask(mask),
        .data_valid(data_mem_valid),
        .valid(instruc_mem_valid),
        .we_re(data_mem_we_re),
        .request(data_mem_request),
        .store_data_out(store_data_out),
        .wrap_load_out(wrap_load_memstage)
    );

    assign rd_memstage = instruction_memstage[11:7];
    assign alu_out_address = alu_res_out_memstage;
    assign mask_singal = mask ;
    assign load_signal = load_memstage;

    //MEMORY STAGE PIPELINE
    memory_pipe u_memstagepipeline(
        .clk(clk),
        .mem_reg_in(mem_to_reg_memstage),
        .wrap_load_in(wrap_load_memstage),
        .alu_res(alu_res_out_memstage),
        .next_sel_addr(next_sel_address_memstage),
        .pre_address_in(pre_pc_addr_memstage),
        .instruction_in(instruction_memstage),
        .reg_write_in(reg_write_memstage),
        .reg_write_out(reg_write_wb),
        .alu_res_out(alu_res_out_wb),
        .mem_reg_out(mem_to_reg_wb),
        .next_sel_address(next_sel_address_wb),
        .instruction_out(instruction_wb),
        .pre_address_out(pre_pc_addr_wb),
        .wrap_load_out(wrap_load_wb)
    );

    //WRITE BACK STAGE
    write_back u_wbstage(
        .mem_to_reg(mem_to_reg_wb),
        .alu_out(alu_res_out_wb),
        .data_mem_out(wrap_load_wb),
        .next_sel_address(next_sel_address_wb),
        .rd_sel_mux_out(rd_wb_data)
    );
endmodule